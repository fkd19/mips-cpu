`timescale 1ns / 1ps

module LED_drive(input LED_WE,
			  input 
    );


endmodule
